interface mux_intf;

logic s;
logic [2:0]a,b;
logic [2:0]y;


modport dut(input a,b,s, output y);


endinterface
